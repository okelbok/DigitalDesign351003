----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 12.02.2026 23:26:29
-- Design Name: 
-- Module Name: or6_gate_primitive - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity OR6 is
port (A, B, C, D, E, F: in std_logic; G: out std_logic);
end OR6;

architecture Behavioral of OR6 is
signal AB, CD, EF, ABCD: std_logic;
begin
AB <= A or B;
CD <= C or D;
ABCD <= AB or CD;
EF <= E or F;
G <= ABCD or EF;
end Behavioral;
